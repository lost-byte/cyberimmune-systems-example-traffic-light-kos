/* Компонент`CSTimes` установка времён переключения режимов */

component traffic_light.CCSMode

endpoints {
    /* именная реализация интерфейса ICSTimes */
    csmode : traffic_light.ICSMode
}
